module
  input    clk,
  input    rst,
  input    int1,
  input    int2,
  input    int3,
  output   out1,
  output   out2,

















endmodule
